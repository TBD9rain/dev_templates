//==================================================================================================
//
//  Project         :
//  File            :
//  Version         :   v0.0.0
//  Title           :
//
//  Description     :
//
//  Additional info :
//  Version history :
//
//  Author          :
//  Email           :
//
//==================================================================================================

module module_name(
    //  IO PORT DECLARATIONS

);

//=======================
//  PARAMETER DEFINITIONS
//=======================



//======================
//  VARIABLE DEFINITIONS
//======================



//===============
//  DESIGN CODING
//===============



endmodule
